//
module top (
);

    system system_i ();
    
endmodule
    
